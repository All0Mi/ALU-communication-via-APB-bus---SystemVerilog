`ifndef ALU_DEF

`define ALU_DEF
`include "./MODEL/apb_exe_unit_3/exe_unit_3/bit_set/bit_set.sv"
`include "./MODEL/apb_exe_unit_3/exe_unit_3/bit_shift/bit_shift.sv"
`include "./MODEL/apb_exe_unit_3/exe_unit_3/comparator/comparator.sv"
`include "./MODEL/apb_exe_unit_3/exe_unit_3/u2_to_sm/u2_to_sm.sv"
`include "./MODEL/apb_exe_unit_3/exe_unit_3/MUX.sv"
`include "./MODEL/apb_exe_unit_3/exe_unit_3/reg.sv"
  
`endif